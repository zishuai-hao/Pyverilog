module top(
    input wire a,    // 输入信号
    output reg out   // 输出信号
);

assign out = 1'b0;
endmodule